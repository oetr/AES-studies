-------------------------------------------------------------------------------
-- Doc: A naive implementation of advanced encryption standard
-------------------------------------------------------------------------------
-- Author    : Peter Samarin <peter.samarin@gmail.com>
-------------------------------------------------------------------------------
-- Copyright (c) 2020 Peter Samarin
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
------------------------------------------------------------
entity AES_Naive is
  port (
    clk              : in    std_logic;
    rst              : in    std_logic);
end entity AES_Naive;
------------------------------------------------------------
architecture arch of AES_Naive is
begin
  
end architecture arch;
